package some_pkg;

	`include "uvm_macros.svh"

	import uvm_pkg::*;

    `include "some_env.sv"
    `include "test_class.sv"

endpackage : some_pkg
